module OR(x, y, out);

input [31:0] x,y;
output [31:0] out;

assign out = a | b;

endmodule